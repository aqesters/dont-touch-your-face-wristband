.title KiCad schematic
U1 SCL +3V3 +3V3 SDA Net-_C2-Pad1_ GND NC_01 GND +3V3 +3V3 INTA2 NC_02 LSM303AGR
C2 Net-_C2-Pad1_ GND 220n
R8 +3V3 Vib+ 22
C7 +3V3 GND 100n
Q1 PB4 GND Vib- 2N7002
TH1 BATT_PRESENT GND 10k therm
R11 Net-_R11-Pad1_ GND 22k
U6 PWR_ON GND PWR_ON NC_03 +3V3 AP2112K-3.3
C9 +BATT GND 4.7u
U4 VDD VDD ~CHRG ~FULL GND Net-_R11-Pad1_ Net-_R12-Pad2_ Net-_R6-Pad1_ +BATT +BATT GND MCP73834
U5 ~RESET INTA2 PB4 GND SDA PB1 SCL +3V3 ATtiny85-20SU
R9 SDA +3V3 4.7k
R10 SCL +3V3 4.7k
R6 Net-_R6-Pad1_ BATT_PRESENT 909
R5 BATT_PRESENT GND 130k
C13 VDD GND 10u
J1 GND VDD Net-_D4-Pad1_ Net-_J1-PadA6_ Net-_J1-PadA7_ NC_04 VDD GND GND VDD Net-_D3-Pad1_ Net-_J1-PadA7_ Net-_J1-PadA6_ NC_05 VDD GND GND USB_C_Receptacle_GCT_USB4085
J2 Vib+ Vib- Conn_01x02_Female
J3 +BATT -BATT Conn_01x02_Female
C11 PWR_ON GND 100n
U2 NC_06 SDA SCL NC_07 GND -BATT ~RESET Net-_R3-Pad1_ +3V3 PWR_ON STC3115AIQT
R3 Net-_R3-Pad1_ BATT_PRESENT 1k
R4 PWR_ON BATT_PRESENT 1M
R2 -BATT GND 50m
R1 +BATT Net-_D1-Pad1_ 220
R14 Net-_D3-Pad1_ GND 5.1k
R13 Net-_D4-Pad1_ GND 5.1k
C12 +3V3 GND 100n
C10 +3V3 GND 100n
C6 +3V3 GND 100n
C4 PWR_ON GND 1u
C5 +3V3 GND 100n
C8 VDD GND 100n
R12 VDD Net-_R12-Pad2_ 1M
D1 Net-_D1-Pad1_ ~CHRG ~FULL PB1 LED_ABGR
C3 +3V3 GND 100n
U3 +3V3 SDA NC_08 SCL +3V3 NC_09 NC_10 GND GND NC_11 VCNL4020-GS08
C1 +3V3 GND 100n
SW1 NC_12 PWR_ON +BATT SW_SPDT
C14 +3V3 GND 47u
D2 VDD GND ESD9B5.0ST5G
D3 Net-_D3-Pad1_ GND ESD9B3.3ST5G
D4 Net-_D4-Pad1_ GND ESD9B3.3ST5G
.end
